library IEEE;
use IEEE.std_logic_1164.all;

entity xnor_gate is
    port(A: in std_logic;     
         B: in std_logic;     
         Y: out std_logic); 
end xnor_gate;

architecture xnorArch of xnor_gate is
 begin
    Y <= (A and B) or (not A and not B)
end xnorArch;
